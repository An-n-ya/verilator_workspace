module example;
    initial begin $display("Hello World4"); $finish; end
endmodule
